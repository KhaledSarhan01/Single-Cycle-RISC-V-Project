module ALU(
    input [31:0] SrcA,
    input [31:0] SrcB,
    output zero,
    output [31:0] ALU_result  
);
 //module behaviour
 /*
 ALU Decoder description is added with the folder 
 zero: it's equal one when ALU_result=0;
 */   
endmodule